package pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;

  `include "xtn.sv"
  `include "agent_config.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "sequencer.sv"
  `include "apb_cov.sv"
  `include "agent.sv"
  `include "seqs.sv"
  
  `include "sbd.sv"
  `include "env.sv"
  `include "test.sv"
endpackage
